fpga_test_project_pll_inst: fpga_test_project_pll
port map(
          REFERENCECLK => ,
          PLLOUTCORE => ,
          PLLOUTGLOBAL => ,
          RESET => 
        );
